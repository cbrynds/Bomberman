module life_bar (
    //ports
);
    
endmodule