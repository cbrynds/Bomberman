module binary_to_bcd (
    input clk, reset, start,
    input [13:0] in,
    output [3:0] bcd3, bcd2, bcd1, bcd0, count,
    output [1:0] state;
); 
    
endmodule